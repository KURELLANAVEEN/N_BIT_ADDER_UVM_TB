package global_values_pkg;
 parameter int N = 4;
endpackage