import uvm_pkg::*; 
`include "uvm_macros.svh"

`include "adder_tb_pkg.sv"
import global_values_pkg::*;

`include "adder_interface.sv"
`include "tb_top.sv"
`include "adder_transaction_item.sv"
`include "adder_sequencer.sv"
`include "adder_driver.sv"
`include "adder_monitor.sv"
`include "adder_agent.sv"
`include "adder_scoreboard.sv"
`include "adder_env.sv"
`include "adder_sequence.sv"
`include "adder_base_test.sv"