package adder_tb_pkg;
  parameter int N = 4;

  `include "adder_transaction_item.sv"
  `include "adder_driver.sv"
endpackage